***** Spice Netlist for Cell 'inverter_tb' *****

************** Module inverter_tb **************
.subckt inverter_tb out in
m0 out in gnd gnd scmosn w='0.6u' l='0.4u' m='1' 
m1 out in vdd vdd scmosp w='1.8u' l='0.4u' m='1' 
.ends inverter_tb
